`timescale 1ns / 1ps

module Execute(

  );

endmodule
