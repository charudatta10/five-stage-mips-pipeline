`timescale 1ns / 1ps

module TestBench();


  initial begin

    #1 $display("Hello, World!");
  end
endmodule
