`timescale 1ns / 1ps

module InstructionFetch(

  );

endmodule
