`timescale 1ns / 1ps

module TestBench();

endmodule
