`timescale 1ns / 1ps

module InstructionDecode(

  );

endmodule
