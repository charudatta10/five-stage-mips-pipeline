`timescale 1ns / 1ps

module WriteBack(

  );

endmodule
